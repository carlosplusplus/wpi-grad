library verilog;
use verilog.vl_types.all;
entity DataPathTester is
end DataPathTester;
