library verilog;
use verilog.vl_types.all;
entity DFlipFlopTester is
end DFlipFlopTester;
