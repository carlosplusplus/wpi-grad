library verilog;
use verilog.vl_types.all;
entity VotingMachineTester is
end VotingMachineTester;
