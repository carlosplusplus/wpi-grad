library verilog;
use verilog.vl_types.all;
entity CompArch_CPU_Tester is
end CompArch_CPU_Tester;
