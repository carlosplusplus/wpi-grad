library verilog;
use verilog.vl_types.all;
entity MemoryModelTester is
end MemoryModelTester;
