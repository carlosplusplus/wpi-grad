library verilog;
use verilog.vl_types.all;
entity FullAdderTester is
end FullAdderTester;
