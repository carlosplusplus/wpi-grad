library verilog;
use verilog.vl_types.all;
entity MooreSeqDetectorTester is
    generic(
        MAX             : integer := 4
    );
end MooreSeqDetectorTester;
