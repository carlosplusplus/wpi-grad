// Carlos Lazo
// ECE574
// Homework #4

// Part 1: Binary Counter, 8bit Implementation
//         using generate statements.

`timescale 1ns/100ps

module BinaryCounter8bit (clk, rst, init, cin, cout);
  
  // Define a parameter so that the adder can be any size:
  
  parameter SIZE = 8;
  
  // Define inputs and outputs:
  
  input  clk, rst, init, cin;
  output cout;
  
  // Variable for moving current cout to the cin of the next adder.
  
  wire   [SIZE-1:0] carry;
  
  genvar i; // Loop variable.
  
  // Generate all instances of counter cells, and link them together.
  
  generate
    
    for (i=0; i < SIZE; i=i+1) begin : counter_cells
      
      // If this is the first run, take in the first
      // cin value, and begin processing accordingly.
      
      if (i == 0)
        CounterCell cc (clk, rst, init, cin, carry[0]);
        
      // If we are at the last index, do the final calculation
      // and set the final carry out value to co.
      
      else if (i == SIZE-1)
        CounterCell cc (clk, rst, init, carry[i-1], cout);
      
      // Otherwise, the current cin is the previous cout,
      // and the current cout is the newly generated cout.
      
      else
        CounterCell cc (clk, rst, init, carry[i-1], carry[i]);
                
    end
 
  endgenerate
  
endmodule