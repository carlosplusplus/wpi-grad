library verilog;
use verilog.vl_types.all;
entity aluCPUTester is
end aluCPUTester;
