library verilog;
use verilog.vl_types.all;
entity minMemValueTester is
end minMemValueTester;
