library verilog;
use verilog.vl_types.all;
entity TextIO is
end TextIO;
