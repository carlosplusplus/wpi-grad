library verilog;
use verilog.vl_types.all;
entity S2PC_Tester is
end S2PC_Tester;
