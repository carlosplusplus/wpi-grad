library verilog;
use verilog.vl_types.all;
entity multTester is
end multTester;
