library verilog;
use verilog.vl_types.all;
entity HW2Pt1Tester is
end HW2Pt1Tester;
