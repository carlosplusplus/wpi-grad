library verilog;
use verilog.vl_types.all;
entity P2SC_Tester is
end P2SC_Tester;
