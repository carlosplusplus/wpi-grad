library verilog;
use verilog.vl_types.all;
entity MealyAndMoore1101Tester is
end MealyAndMoore1101Tester;
