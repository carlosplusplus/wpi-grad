library verilog;
use verilog.vl_types.all;
entity P2SC_To_S2PC_Tester is
end P2SC_To_S2PC_Tester;
