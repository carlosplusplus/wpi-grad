library verilog;
use verilog.vl_types.all;
entity BoothMultiplier_Testbench is
end BoothMultiplier_Testbench;
