library verilog;
use verilog.vl_types.all;
entity S2PC_To_P2SC_Tester is
end S2PC_To_P2SC_Tester;
