library verilog;
use verilog.vl_types.all;
entity MooreDetector1101Tester is
end MooreDetector1101Tester;
