library verilog;
use verilog.vl_types.all;
entity transistorCircuitTestbench is
end transistorCircuitTestbench;
