library verilog;
use verilog.vl_types.all;
entity ALU16bitModelComparison is
    generic(
        SIM_CHOICE      : integer := 5
    );
end ALU16bitModelComparison;
