library verilog;
use verilog.vl_types.all;
entity FullAdder4bit_Pt3Tester is
    generic(
        SIZE            : integer := 4;
        SIM_CHOICE      : integer := 2
    );
end FullAdder4bit_Pt3Tester;
