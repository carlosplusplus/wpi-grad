library verilog;
use verilog.vl_types.all;
entity ALU16bitTimeTest is
end ALU16bitTimeTest;
