library verilog;
use verilog.vl_types.all;
entity rtlRouterTester is
end rtlRouterTester;
