library verilog;
use verilog.vl_types.all;
entity BinaryCounter8bitTester is
    generic(
        SIZE            : integer := 8
    );
end BinaryCounter8bitTester;
