library verilog;
use verilog.vl_types.all;
entity ALU2bitTester is
end ALU2bitTester;
