library verilog;
use verilog.vl_types.all;
entity ALU8bitTester is
end ALU8bitTester;
